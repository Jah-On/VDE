module vlang

import gx 

pub const (
	kw_map = {
		"as":        gx.rgb(180, 0, 180)
		"asm":       gx.rgb(220, 0, 220)
		"assert":    gx.rgb(220, 0, 220)
		"atomic":    gx.rgb(0, 255, 25)
		"break":     gx.rgb(220, 0, 220)
		"const":     gx.rgb(220, 0, 220)
		"continue":  gx.rgb(220, 0, 220)
		"defer":     gx.rgb(220, 0, 220)
		"dump":      gx.rgb(150, 0, 0)
		"else":      gx.rgb(220, 0, 220)
		"enum":      gx.rgb(120, 120, 120)
		"false":     gx.rgb(0, 0, 255)
		"for":       gx.rgb(220, 0, 220)
		"fn":        gx.rgb(255, 255, 128)
		"global":    gx.rgb(220, 0, 220)
		"go":        gx.rgb(220, 0, 220)
		"goto":      gx.rgb(220, 0, 220)
		"if":        gx.rgb(220, 0, 220)
		"import":    gx.rgb(180, 0, 180)
		"in":        gx.rgb(220, 0, 220)
		"interface": gx.rgb(140, 0, 140)
		"is":        gx.rgb(220, 0, 220)
		"lock":      gx.rgb(220, 0, 220)
		"match":     gx.rgb(220, 0, 220)
		"module":    gx.rgb(180, 0, 180)
		"mut":       gx.rgb(255, 200, 0)
		"none":      gx.rgb(100, 0, 0)
		"offsetof":  gx.rgb(150, 0, 0)
		"orelse":    gx.rgb(220, 0, 220)
		"pub":       gx.rgb(255, 200, 0)
		"rlock":     gx.rgb(220, 0, 220)
		"select":    gx.rgb(220, 0, 220)
		"sizeof":    gx.rgb(150, 0, 0)
		"shared":    gx.rgb(255, 200, 0)
		"static":    gx.rgb(255, 200, 0)
		"struct":    gx.rgb(100, 100, 100)
		"true":      gx.rgb(0, 0, 255)
		"type":      gx.rgb(180, 180, 180)
		"typeof":    gx.rgb(150, 0, 0)
		"union":     gx.rgb(160, 160, 160)
		"unsafe":    gx.rgb(220, 0, 220)
		"bool":      gx.rgb(0, 0, 255)
		"i8":        gx.rgb(50, 100, 255)
		"i16":       gx.rgb(50, 100, 255)
		"int":       gx.rgb(50, 100, 255)
		"i64":       gx.rgb(50, 100, 255)
		"u8":        gx.rgb(50, 150, 255)
		"u16":       gx.rgb(50, 150, 255)
		"u32":       gx.rgb(50, 150, 255)
		"u64":       gx.rgb(50, 150, 255)
		"f32":       gx.rgb(0, 200, 255)
		"f64":       gx.rgb(0, 200, 255)
		"string":    gx.rgb(0, 200, 100)
		"rune":      gx.rgb(0, 150, 50)
		"voidptr":   gx.rgb(100, 0, 0)
	}
	kw_list = kw_map.keys()
)